///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Standard Covergroups
//
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file
// except in compliance with the License, or, at your option, the Apache License version 2.0. You
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,
// either express or implied. See the License for the specific language governing permissions
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////

`define RAMBASEADDR 32'h80000000
`define LARGESTPROGRAM 32'h00010000
`define SAFEREGIONSTART (`RAMBASEADDR + `LARGESTPROGRAM)
`define REGIONSTART `SAFEREGIONSTART

`define COVER_RV32PMP
`define COVER_RV64PMP

covergroup PMPM_cfg0_cg with function sample(ins_t ins);
    option.per_instance = 0;
    `include  "coverage/RISCV_coverage_standard_coverpoints.svh"

    rs1_in_region: coverpoint ins.current.rs1_val {
        bins at_region     = {`REGIONSTART};
    }

    Mcause: coverpoint ins.current.csr[12'h342]{  
        bins illegal_ins  = {32'd2};
        bins no_exception = {32'd0};
    }

    exec_instr: coverpoint ins.current.insn {
        wildcard bins jalr = {32'b????????????_?????_000_?????_1100111};
    }

    read_instr: coverpoint ins.current.insn {
        wildcard bins lb  = {32'b????????????_?????_000_?????_0000011};
        wildcard bins lbu = {32'b????????????_?????_100_?????_0000011};
        wildcard bins lh  = {32'b????????????_?????_001_?????_0000011};
        wildcard bins lhu = {32'b????????????_?????_101_?????_0000011};
        wildcard bins lw  = {32'b????????????_?????_010_?????_0000011};
        `ifdef XLEN64
            wildcard bins lwu = {32'b????????????_?????_110_?????_0000011};
            wildcard bins ld  = {32'b????????????_?????_011_?????_0000011};
        `endif
    }

    write_instr: coverpoint ins.current.insn {
        wildcard bins sb = {32'b?????????_?????_?????_000_?????_0100011};
        wildcard bins sh = {32'b?????????_?????_?????_001_?????_0100011};
        wildcard bins sw = {32'b?????????_?????_?????_010_?????_0100011};
        `ifdef XLEN64
            wildcard bins sd = {32'b?????????_?????_?????_011_?????_0100011};
        `endif
    }

    fetch_result: coverpoint ins.current.csr[12'h342] { 
        bins instr_access_fault = {32'd1};
        bins no_exception = {32'd0};
    }

    read_result: coverpoint ins.current.csr[12'h342] { 
        bins load_access_fault = {32'd5};
        bins no_exception = {32'd0};
    }

    write_result: coverpoint ins.current.csr[12'h342] { 
        bins store_access_fault = {32'd7};
        bins no_exception = {32'd0};
    }

    legal_lxwr_cfg0: coverpoint ins.current.csr[12'h3A0][7:0] { // For both RV32 and RV64
        wildcard bins cfg_l000 = {8'b10011000};
        wildcard bins cfg_l001 = {8'b10011001};
        wildcard bins cfg_l011 = {8'b10011011};
        wildcard bins cfg_l100 = {8'b10011100};
        wildcard bins cfg_l101 = {8'b10011101};
        wildcard bins cfg_l111 = {8'b10011111};
    }

    pmpcfg0_L0_all: coverpoint ins.current.csr[12'h3A0] {
        `ifdef XLEN32
            wildcard bins pmp0cfg_L0  = {32'b????????????????????????00011000};
            wildcard bins pmp1cfg_L0  = {32'b????????????????00011000????????};
            wildcard bins pmp2cfg_L0  = {32'b????????00011000????????????????};
            wildcard bins pmp3cfg_L0  = {32'b00011000????????????????????????};
        `endif
        `ifdef XLEN64
            wildcard bins pmp0cfg_L0  = {64'b????????????????????????????????????????????????????????00011000};
            wildcard bins pmp1cfg_L0  = {64'b????????????????????????????????????????00011000????????????????};
            wildcard bins pmp2cfg_L0  = {64'b????????????????????????00011000????????????????????????????????};
            wildcard bins pmp3cfg_L0  = {64'b????????00011000????????????????????????????????????????????????};
        `endif
    }

    pmpcfg0_X0_all: coverpoint ins.current.csr[12'h3A0] {
        `ifdef XLEN32
            wildcard bins pmp0cfg_X0  = {32'b????????????????????????100110??};
            wildcard bins pmp1cfg_X0  = {32'b????????????????100110??????????};
            wildcard bins pmp2cfg_X0  = {32'b????????100110??????????????????};
            wildcard bins pmp3cfg_X0  = {32'b100110??????????????????????????};
        `endif
        `ifdef XLEN64
            wildcard bins pmp0cfg_X0  = {64'b????????????????????????????????????????????????????????100110??};
            wildcard bins pmp1cfg_X0  = {64'b????????????????????????????????????????100110??????????????????};
            wildcard bins pmp2cfg_X0  = {64'b????????????????????????100110??????????????????????????????????};
            wildcard bins pmp3cfg_X0  = {64'b????????100110??????????????????????????????????????????????????};
        `endif
    }

    pmpcfg0_X1_all: coverpoint ins.current.csr[12'h3A0] {
        `ifdef XLEN32
            wildcard bins pmp0cfg_X1  = {32'b????????????????????????100111??};
            wildcard bins pmp1cfg_X1  = {32'b????????????????100111??????????};
            wildcard bins pmp2cfg_X1  = {32'b????????100111??????????????????};
            wildcard bins pmp3cfg_X1  = {32'b100111??????????????????????????};
        `endif
        `ifdef XLEN64
            wildcard bins pmp0cfg_X1  = {64'b????????????????????????????????????????????????????????100111??};
            wildcard bins pmp1cfg_X1  = {64'b????????????????????????????????????????100111??????????????????};
            wildcard bins pmp2cfg_X1  = {64'b????????????????????????100111??????????????????????????????????};
            wildcard bins pmp3cfg_X1  = {64'b????????100111??????????????????????????????????????????????????};
        `endif
    }

    pmpcfg0_RW00_all: coverpoint ins.current.csr[12'h3A0] {
        `ifdef XLEN32
            wildcard bins pmp0cfg_RW00  = {32'b????????????????????????10011100};
            wildcard bins pmp1cfg_RW00  = {32'b????????????????10011100????????};
            wildcard bins pmp2cfg_RW00  = {32'b????????10011100????????????????};
            wildcard bins pmp3cfg_RW00  = {32'b10011100????????????????????????};
        `endif
        `ifdef XLEN64
            wildcard bins pmp0cfg_RW00  = {64'b????????????????????????????????????????????????????????10011100};
            wildcard bins pmp1cfg_RW00  = {64'b????????????????????????????????????????10011100????????????????};
            wildcard bins pmp2cfg_RW00  = {64'b????????????????????????10011100????????????????????????????????};
            wildcard bins pmp3cfg_RW00  = {64'b????????10011100????????????????????????????????????????????????};
        `endif
    }

    pmpcfg0_RW10_all: coverpoint ins.current.csr[12'h3A0] {
        `ifdef XLEN32
            wildcard bins pmp0cfg_RW10  = {32'b????????????????????????10011101};
            wildcard bins pmp1cfg_RW10  = {32'b????????????????10011101????????};
            wildcard bins pmp2cfg_RW10  = {32'b????????10011101????????????????};
            wildcard bins pmp3cfg_RW10  = {32'b10011101????????????????????????};
        `endif
        `ifdef XLEN64
            wildcard bins pmp0cfg_RW10  = {64'b????????????????????????????????????????????????????????10011101};
            wildcard bins pmp1cfg_RW10  = {64'b????????????????????????????????????????10011101????????????????};
            wildcard bins pmp2cfg_RW10  = {64'b????????????????????????10011101????????????????????????????????};
            wildcard bins pmp3cfg_RW10  = {64'b????????10011101????????????????????????????????????????????????};
        `endif
    }

    pmpcfg0_RW11_all: coverpoint ins.current.csr[12'h3A0] {
        `ifdef XLEN32
            wildcard bins pmp0cfg_RW11  = {32'b????????????????????????10011111};
            wildcard bins pmp1cfg_RW11  = {32'b????????????????10011111????????};
            wildcard bins pmp2cfg_RW11  = {32'b????????10011111????????????????};
            wildcard bins pmp3cfg_RW11  = {32'b10011111????????????????????????};
        `endif
        `ifdef XLEN64
            wildcard bins pmp0cfg_RW11  = {64'b????????????????????????????????????????????????????????10011111};
            wildcard bins pmp1cfg_RW11  = {64'b????????????????????????????????????????10011111????????????????};
            wildcard bins pmp2cfg_RW11  = {64'b????????????????????????10011111????????????????????????????????};
            wildcard bins pmp3cfg_RW11  = {64'b????????10011111????????????????????????????????????????????????};
        `endif
    }

    cp_cfg_X_set: cross legal_lxwr_cfg0, fetch_result, exec_instr, rs1_in_region {
        ignore_bins ig1 = binsof(legal_lxwr_cfg0.cfg_l000);
        ignore_bins ig2 = binsof(legal_lxwr_cfg0.cfg_l001);
        ignore_bins ig3 = binsof(legal_lxwr_cfg0.cfg_l011);
        ignore_bins ig4 = binsof(fetch_result.instr_access_fault);
    }

    cp_cfg_X_unset: cross legal_lxwr_cfg0, fetch_result, exec_instr, rs1_in_region {
        ignore_bins ig1 = binsof(legal_lxwr_cfg0.cfg_l100);
        ignore_bins ig2 = binsof(legal_lxwr_cfg0.cfg_l101);
        ignore_bins ig3 = binsof(legal_lxwr_cfg0.cfg_l111);
        ignore_bins ig4 = binsof(fetch_result.no_exception);
    }

    cp_cfg_R_set: cross legal_lxwr_cfg0, read_result, read_instr, rs1_in_region {
        ignore_bins ig1 = binsof(legal_lxwr_cfg0.cfg_l000);
        ignore_bins ig2 = binsof(legal_lxwr_cfg0.cfg_l100);
        ignore_bins ig3 = binsof(read_result.load_access_fault);
    }

    cp_cfg_R_unset: cross legal_lxwr_cfg0, read_result, read_instr, rs1_in_region {
        ignore_bins ig1 = binsof(legal_lxwr_cfg0.cfg_l001);
        ignore_bins ig2 = binsof(legal_lxwr_cfg0.cfg_l011);
        ignore_bins ig3 = binsof(legal_lxwr_cfg0.cfg_l101);
        ignore_bins ig4 = binsof(legal_lxwr_cfg0.cfg_l111);
        ignore_bins ig5 = binsof(read_result.no_exception);
    }

    cp_cfg_W_set: cross legal_lxwr_cfg0, write_result, write_instr, rs1_in_region {
        ignore_bins ig1 = binsof(legal_lxwr_cfg0.cfg_l000);
        ignore_bins ig2 = binsof(legal_lxwr_cfg0.cfg_l001);
        ignore_bins ig3 = binsof(legal_lxwr_cfg0.cfg_l101);
        ignore_bins ig4 = binsof(legal_lxwr_cfg0.cfg_l100);
        ignore_bins ig5 = binsof(write_result.store_access_fault);
    }

    cp_cfg_W_unset: cross legal_lxwr_cfg0, write_result, write_instr, rs1_in_region {
        ignore_bins ig1 = binsof(legal_lxwr_cfg0.cfg_l011);
        ignore_bins ig2 = binsof(legal_lxwr_cfg0.cfg_l111);
        ignore_bins ig3 = binsof(write_result.no_exception);
    }

    cp_cfg_X0_all: cross pmpcfg0_X0_all, fetch_result, exec_instr, rs1_in_region {  // For first four regions.
        ignore_bins ig1 = binsof(fetch_result.no_exception);
    }

    cp_cfg_X1_all: cross pmpcfg0_X1_all, fetch_result, exec_instr, rs1_in_region { // For first four regions.
        ignore_bins ig1 = binsof(fetch_result.instr_access_fault);
    }

    cp_cfg_RW00_all: cross pmpcfg0_RW00_all, read_result, write_result, rs1_in_region { // For first four regions.
        ignore_bins ig1 = binsof(read_result.no_exception);
        ignore_bins ig2 = binsof(write_result.no_exception);
    }

    cp_cfg_RW10_all: cross pmpcfg0_RW10_all, read_result, write_result, rs1_in_region { // For first four regions.
        ignore_bins ig1 = binsof(read_result.load_access_fault);
        ignore_bins ig2 = binsof(write_result.no_exception);
    }

    cp_cfg_RW11_all: cross pmpcfg0_RW11_all, read_result, write_result, rs1_in_region { // For first four regions.
        ignore_bins ig1 = binsof(read_result.load_access_fault);
        ignore_bins ig2 = binsof(write_result.store_access_fault);
    }
    
    cp_cfg_L_access_all: cross pmpcfg0_L0_all, exec_instr, read_instr, write_instr, Mcause, rs1_in_region { // For first four regions.
        ignore_bins ig1 = binsof(Mcause.illegal_ins);
        ignore_bins ig2 = binsof(read_instr.lh);
        ignore_bins ig3 = binsof(read_instr.lhu);
        ignore_bins ig4 = binsof(read_instr.lb);
        ignore_bins ig5 = binsof(read_instr.lbu);
        ignore_bins ig6 = binsof(write_instr.sh);
        ignore_bins ig7 = binsof(write_instr.sb);
        `ifdef XLEN64
            ignore_bins ig8 = binsof(read_instr.lwu);
            ignore_bins ig9 = binsof(read_instr.ld);
            ignore_bins ig10 = binsof(write_instr.sd);
        `endif
    } 
 
endgroup

function void pmp_sample(int hart, int issue, ins_t ins);
    PMPM_cfg0_cg.sample(ins);
endfunction
